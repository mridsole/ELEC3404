*** ELEC3404 Lab 2 Amplifier Circuit ***

R1 VCC B 27k
R2 B GND 150k
RC VCC C 8.2k
RE E GND 1.8k

Q1 C B E BC547

* voltage source:
VS VCC GND DC 20 AC 0

* https://github.com/saketkc/kicad-ngspice/blob/master/modelEditor_mail/BC547.txt
.model BC547 NPN( Vtf=1.7 Cjc=7.306p Nc=2 Tr=46.91n Ne=1.307 
+ Cje=22.01p Isc=0 Xtb=1.5 Rb=10 Rc=1 
+ Tf=411.1p Xti=3 Ikr=0 Bf=213 Fc=.5 
+ Ise=14.34f Br=6.092 Ikf=.2847 Mje=.377 Mjc=.3416 
+ Vaf=74.03 Vjc=.75 Vje=.75 Xtf=3 Itf=.6 
+ Is=14.34f Eg=1.11 )

.end
