.model 1N914 D(Is=2.52n Rs=0.568 N=1.752 Cjo=4p M=.4 tt=20n Iave=200m Vpk=75 mfg=Motorola type=silicon )
.model 1N4148 D(Is=2.52n Rs=0.568 N=1.752 Cjo=4p M=.4 tt=20n Iave=200m Vpk=75 mfg=Motorola type=silicon )
.model MMSD4148 D(Is=2.52n Rs=0.568 N=1.752 Cjo=.64p M=.4 tt=5n Iave=200m Vpk=100 mfg=Onsemi type=silicon )
.model 1N5817 D(Is=31.7u Rs=0.051 N=1.373 Cjo=190p M=.3 Eg=.69 Xti=2 Iave=1 Vpk=20 mfg=Motorola type=Schottky)
.model 1N5818 D(Is=31.7u Rs=0.051 N=1.373 Cjo=160p M=.38 Eg=.69 Xti=2 Iave=1 Vpk=30 mfg=Motorola type=Schottky)
.model 1N5819 D(Is=31.7u Rs=0.051 N=1.373 Cjo=110p M=.35 Eg=.69 Xti=2 Iave=1 Vpk=40 mfg=Motorola type=Schottky)
.model BAT54 D(Is=.1u Rs=2.2 N=1 Cjo=12p M=.3 Eg=.69 Xti=2 Iave=300m Vpk=30 mfg=Vishay type=Schottky)
.model MBR0520L D(Is=82.5n Rs=0.115 N=.7228 Cjo=180p M=.63 Eg=.69 Xti=2 Iave=.5 Vpk=20 mfg=Motorola type=Schottky)
.model MBR0530L D(Is=1.55u Rs=0.0858 N=1.079 Cjo=180p Eg=.69 Xti=2 Iave=.5 Vpk=30 mfg=Motorola type=Schottky)
.model MBRS1100 D(Is=20.6u Rs=0.0079 N=2.303 Cjo=270p M=.575 Eg=.69 Xti=2 Iave=1 Vpk=100 mfg=Motorola type=Schottky)
.model MBRS130L D(Is=772n Rs=0.0299 N=.8442 Cjo=290p M=.7 Eg=.69 Xti=2 Iave=1 Vpk=30 mfg=Motorola type=Schottky)
.model MBRS140 D(Is=235n Rs=0.109 N=.7760 Cjo=160p M=.6 Eg=.69 Xti=2 Iave=1 Vpk=40 mfg=Motorola type=Schottky)
.model MBRS340 D(Is=22.6u Rs=0.042 N=1.094 Cjo=480p M=.61 Eg=.69 Xti=2 Iave=3 Vpk=40 mfg=Motorola type=Schottky)
.model MBRS360 D(Is=22.6u Rs=0.042 N=1.094 Cjo=480p M=.61 Eg=.69 Xti=2 Iave=3 Vpk=60 mfg=Motorola type=Schottky)
.model CMDSH2-3 D(Is=210nA Rs=0.5 N=1.09 Cjo=50p M=.5 Eg=.69 Xti=2 Iave=200m Vpk=30 mfg=Central type=Schottky)
.model MURS120 D(Is=33.8n Rs=0.0236 N=1.718 Cjo=45p M=.6 tt=45n Iave=1 Vpk=200 mfg=Motorola type=silicon )
.model MURS320 D(Is=1.06n Rs=0.0111 N=1.367 Cjo=135p M=.45 tt=45n Iave=3 Vpk=200 mfg=Motorola type=silicon )
.model MBR735 D(Is=159u Rs=0.02 N=1.76 Cjo=740p M=.6 Eg=.69 Xti=2 Iave=7.5 Vpk=35 mfg=Motorola type=Schottky)
.model MBR745 D(Is=159u Rs=0.02 N=1.76 Cjo=740p M=.6 Eg=.69 Xti=2 Iave=7.5 Vpk=45 mfg=Motorola type=Schottky)
.model BZX84C6V2L D(Is=1.5n Rs=.5 Cjo=185p nbv=3 bv=6.2 Ibv=1m Vpk=6.2 mfg=Motorola type=zener )
.model BZX84C8V2L D(Is=0.8n Rs=.5 Cjo=135p nbv=3 bv=8.2 Ibv=1m Vpk=8.2 mfg=Motorola type=zener )
.model BZX84C10L D(Is=0.6u Rs=.5 Cjo=150p nbv=5 bv=10 Ibv=1m Vpk=10 mfg=Motorola type=zener )
.model BZX84C12L D(Is=0.6u Rs=.5 Cjo=150p nbv=5 bv=12 Ibv=1m Vpk=12 mfg=Motorola type=zener )
.model BZX84C15L D(Is=0.6u Rs=.5 Cjo=110p nbv=6 bv=15 Ibv=1m Vpk=15 mfg=Motorola type=zener )
.model RB10L-40 D(Is=2.6uA Rs=0.0674 N=1.163 Cjo=180p M=.6 Eg=.69 Xti=2 Iave=1 Vpk=40 mfg=Rohm type=Schottky)
.model 1N750 D(Is=.88f Rs=.25 Cjo=175p M=.55 nbv=1.7 bv=4.7 Vj=.75 Isr=1.86n Nr=2 Ibv=20.245m Ibvl=1.96m Nbvl=15 Tbv1=-21.3u Vpk=4.7 mfg=Motorola type=zener)
.model MV2201 D(Is=1.365p Rs=1 Cjo=14.93p M=.4261 Vj=.75 Isr=16.02p Nr=2 Bv=25 Ibv=10u Vpk=25 mfg=Motorola type=varactor)
.model MBR0540 D(Is=9.11u Rs=0.121 N=1.33753 Eg=0.69 Xti=2 Cjo=194p Vj=0.25 M=.4 Iave=.5 Vpk=40 mfg=GI type=Schottky)
.model MUR460 D(Is=149n Rs=0.0384 N=2 EG=1.285 XTI=0.5 BV=800 IBV=1e-05 Cjo=126.4p Vj=1.34 M=0.52 tt=44.4n Iave=4 Vpk=600 mfg=GI type=silicon)
.model MBRB2545CT D(Is=19.4n Rs=0.01 N=0.733 Eg=0.718 Xti=0.535 Cjo=2.05n Vj=0.4 M=0.41 Iave=25 Vpk=45 mfg=GI type=Schottky)
.model MBR20100CT D(Is=10u Rs=0.005 N=1.5 Ikf=.3 Isr=10u Nr=3 Cjo=1e-11 Vj=0.7 Iave=10 Vpk=100 mfg=Motorola type=Schottky)
.model 30BQ060 D(Is=10u Rs=0.04 N=1.4 Cjo=180p Eg=.69 Xti=2 Iave=3 Vpk=60 mfg=International_Rectifier type=Schottky)
.model UPSC600 D(Is=2p Rs=0.33 N=1.5 Cjo=50p M=.3 Iave=1 Vpk=600 mfg=Microsemi type=SiC_Schottky)
.model NSPW500BS D(Is=0.27n Rs=5.65 N=6.79 Cjo=42p Iave=30m Vpk=5 mfg=Nichia type=LED)
.model QTLP690C D(Is=1e-22 Rs=6 N=1.5 Cjo=50p Iave=160m Vpk=5 mfg=Fairchild type=LED)
.model PMEG2020AEA D(Is=5.409u Rs=0.05676 N=1.02 Cjo=0.1908n M=0.4863 Eg=0.69 Xti=2 BV=22 IBV=50u Vj=0.3408 FC=0.5 Iave=2 Vpk=20 mfg=Philips type=Schottky)
.model PMEG2010EA D(Is=1.686u Rs=0.1249 N=1.015 Cjo=90.86p M=0.4542 Eg=0.69 Xti=2 BV=21 IBV=1u Vj=0.1939 FC=1 Iave=1 Vpk=20 mfg=Philips type=Schottky)
.model PMEG2010BEA D(Is=3.334u Rs=0.08222 N=0.9791 Cjo=0.1266n M=0.5 Eg=0.69 Xti=2 BV=22 IBV=0.0001 Vj=0.3619 FC=0.5 Iave=1 Vpk=20 mfg=Philips type=Schottky)
.model PMEG3010BEA D(Is=2.936u Rs=0.1166 N=0.9839 Cjo=0.1068n M=0.4948 Eg=0.69 Xti=2 BV=33 IBV=75u Vj=0.3459 FC=0.5 Iave=1 Vpk=30 mfg=Philips type=Schottky)
.model PMEG4010BEA D(Is=2.831u Rs=0.1975 N=0.9816 Cjo=84.37p M=0.4789 Eg=0.69 Xti=2 BV=44 IBV=50u Vj=0.3116 FC=0.5 Iave=1 Vpk=40 mfg=Philips type=Schottky)
.model PMEG2005AEA D(Is=3.334u Rs=0.08222 N=0.9791 Cjo=0.1266n M=0.5 Eg=0.69 Xti=2 BV=22 IBV=0.0001 Vj=0.3619 FC=0.5 Iave=0.5 Vpk=20 mfg=Philips type=Schottky)
.model PMEG3005AEA D(Is=2.936u Rs=0.1166 N=0.9839 Cjo=0.1068n M=0.4948 Eg=0.69 Xti=2 BV=33 IBV=75u Vj=0.3459 FC=0.5 Iave=0.5 Vpk=30 mfg=Philips type=Schottky)
.model PMEG4005AEA D(Is=2.831u Rs=0.1975 N=0.9816 Cjo=84.37p M=0.4789 Eg=0.69 Xti=2 BV=44 IBV=50u Vj=0.3116 FC=0.5 Iave=0.5 Vpk=40 mfg=Philips type=Schottky)
.model PMEG2010AEB D(Is=87.24u Rs=0.2728 N=0.9699 Cjo=29.99p M=0.3755 Eg=0.69 Xti=2 BV=22 IBV=0.0004 Vj=0.2604 FC=0.5 Iave=1 Vpk=20 mfg=Philips type=Schottky)
.model PMEG2005EB D(Is=0.9985u Rs=0.2146 N=0.9283 Cjo=61.05p M=0.4159 Eg=0.69 Xti=2 BV=32 IBV=0.001 Vj=0.1 FC=0.5 Iave=0.5 Vpk=20 mfg=Philips type=Schottky)
.model PMEG6010AED D(Is=0.5u Rs=0.3422 N=0.9751 Cjo=0.175n M=0.4725 Eg=0.69 Xti=2 BV=66 IBV=0.0004 Vj=0.3761 FC=0.5 Iave=1 Vpk=60 mfg=Philips type=Schottky)
.model PRLL5817 D(Is=2.119u Rs=0.0419 N=1.02 Cjo=0.252n M=0.5104 Eg=0.69 Xti=2 BV=1000 IBV=0.001 Vj=0.4792 FC=0.5 Iave=1 Vpk=20 mfg=Philips type=Schottky)
.model LXHL-BW02 D(Is=4.5e-20 Rs=0.85 N=2.6 Cjo=1.18n Iave=400mA mfg=Lumileds type=LED)
.model GSD2004W-V D(Is=1e-14 Rs=1.6 N=1 Cjo=5p tt=50n Iave=225m Vpk=300 mfg=Vishay type=silicon)
.MODEL IN4007 D(IS=7.02767e-09 RS=0.0341512 N=1.80803 EG=1.05743 XTI=5 BV=1000 IBV=5e-08 CJO=1e-11 VJ=0.7 M=0.5 FC=0.5 TT=1e-07 KF=0 AF=1)
.MODEL D1N4001 D(IS=29.5E-9 RS=73.5E-3 N=1.96 CJO=34.6P VJ=0.627 M=0.461 BV=60 IBV=10U)

.model 2N2222 NPN(IS=1E-14 VAF=100 BF=200 IKF=0.3 XTB=1.5 BR=3 CJC=8E-12 CJE=25E-12 TR=100E-9 TF=400E-12 ITF=1 VTF=2 XTF=3 RB=10 RC=3 RE=1 Vceo=30 Icrating=800m mfg=Philips)
.model 2N2907 PNP(IS=1E-14 VAF=120 BF=250 IKF=0.3 XTB=1.5 BR=3 CJC=8E-12 CJE=30E-12 TR=100E-9 TF=400E-12 ITF=1 VTF=2 XTF=3 RB=10 RC=3 RE=1 Vceo=40 Icrating=600m mfg=Philips)
.model 2N3904 NPN(IS=1E-14 VAF=100 Bf=300 IKF=0.4 XTB=1.5 BR=4 CJC=4E-12 CJE=8E-12 RB=20 RC=0.1 RE=0.1 TR=250E-9 TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m mfg=Philips)
.model 2N3906 PNP(IS=1E-14 VAF=100 BF=200 IKF=0.4 XTB=1.5 BR=4 CJC=4.5E-12 CJE=10E-12 RB=20 RC=0.1 RE=0.1 TR=250E-9 TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m mfg=Philips)
.model FZT849 NPN(IS=5.8591E-13 NF=0.9919 BF=230 IKF=18 VAF=90 ISE=2.0067E-13 NE=1.4 NR=0.9908 BR=180 IKR=6.8 VAR=20 ISC=5.3E-13 NC=1.46 RB=0.023 RE=0.0223 RC=0.015 CJC=200E-12 MJC=0.3006 VJC=0.3532 CJE=1.21E-9 TF=1.07E-9 TR=9.3E-9 Vceo=30 Icrating=7 mfg=Zetex) ; Zetex PLC, Fields New Road, Chadderton, Oldham OL9 8NP
.model ZTX849 ako:FZT849 NPN(Vceo=30 Icrating=7 mfg=Zetex)
.model ZTX1048A NPN(IS=13.73E-13 NF=1.0 BF=550 IKF=8.0 VAF=120 ISE=2.6E-13 NE=1.38 NR=1.0 BR=300 IKR=6 VAR=15 ISC=1.6E-12 NC=1.4 RB=0.1 RE=0.022 RC=0.010 CJC=136E-12 CJE=559.1E-12 MJC=0.267 MJE=0.299 VJC=0.420 VJE=0.533 TF=600E-12 TR=3E-9 Vceo=17.5 Icrating=5 mfg=Zetex) ; Zetex PLC, Fields New Road, Chadderton, Oldham OL9 8NP
.model 2N4124 NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=495 Ne=1.28 Ise=6.734f Ikf=69.35m Xtb=1.5 Br=.7214 Nc=2 Isc=0 Ikr=0 Rc=1 Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75 Tr=238.3n Tf=301.3p Itf=.4 Vtf=4 Xtf=2 Rb=10 Vceo=25 Icrating=200m mfg=Fairchild)
.model 2N4126 PNP(Is=1.41f Xti=3 Eg=1.11 Vaf=18.7 Bf=203.7 Ne=1.5 Ise=0 Ikf=80m Xtb=1.5 Br=4.924 Nc=2 Isc=0 Ikr=0 Rc=2.5 Cjc=9.728p Mjc=.5776 Vjc=.75 Fc=.5 Cje=8.063p Mje=.3677 Vje=.75 Tr=33.23n Tf=179.3p Itf=.4 Vtf=4 Xtf=6 Rb=10 Rb=10 Vceo=25 Icrating=200m mfg=Fairchild)
.model 2N3391A NPN(Is=12.03f Xti=3 Eg=1.11 Vaf=37.37 Bf=427.8 Ne=1.971 Ise=2.953p Ikf=.1072 Xtb=1.5 Br=4.379 Nc=2 Isc=0 Ikr=0 Rc=1 Cjc=5.777p Mjc=.3199 Vjc=.75 Fc=.5 Cje=8.307p Mje=.384 Vje=.75 Tr=701.7p Tf=385.4p Itf=.17 Vtf=3 Xtf=8 Rb=10 Vceo=25 Icrating=500m mfg=Fairchild)
.model 2N5089 NPN(Is=5.911f Xti=3 Eg=1.11 Vaf=62.37 Bf=1.434K Ne=1.421 Ise=5.911f Ikf=15.4m Xtb=1.5 Br=1.262 Nc=2 Isc=0 Ikr=0 Rc=1.61 Cjc=4.017p Mjc=.3174 Vjc=.75 Fc=.5 Cje=4.973p Mje=.4146 Vje=.75 Tr=4.671n Tf=822.3p Itf=.35 Vtf=4 Xtf=7 Rb=10 Vceo=25 Icrating=100m mfg=Fairchild)
.model 2N5210 NPN(Is=5.911f Xti=3 Eg=1.11 Vaf=62.37 Bf=809.9 Ne=1.358 Ise=5.911f Ikf=14.26m Xtb=1.5 Br=1.287 Nc=2 Isc=0 Ikr=0 Rc=1.61 Cjc=4.017p Mjc=.3174 Vjc=.75 Fc=.5 Cje=4.973p Mje=.4146 Vje=.75 Tr=4.68n Tf=820.9p Itf=.35 Vtf=4 Xtf=7 Rb=10 Vceo=50 Icrating=100m mfg=Fairchild)
.model 2N5087 PNP(Is=6.734f Xti=3 Eg=1.11 Vaf=45.7 Bf=254.1 Ne=1.741 Ise=6.734f Ikf=.1962 Xtb=1.5 Br=2.683 Nc=2 Isc=0 Ikr=0 Rc=1.67 Cjc=6.2p Mjc=.301 Vjc=.75 Fc=.5 Cje=7.5p Mje=.2861 Vje=.75 Tr=10.1n Tf=467.8p Itf=.17 Vtf=5 Xtf=8 Rb=10 Vceo=50 Icrating=100m mfg=Fairchild)
.model 2N2219A NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=74.03 Bf=255.9 Ne=1.307 Ise=14.34f Ikf=.2847 Xtb=1.5 Br=6.092 Nc=2 Isc=0 Ikr=0 Rc=1 Cjc=7.306p Mjc=.3416 Vjc=.75 Fc=.5 Cje=22.01p Mje=.377 Vje=.75 Tr=46.91n Tf=411.1p Itf=.6 Vtf=1.7 Xtf=3 Rb=10 Vceo=40 Icrating=800m mfg=Philips)
.model 2N2905A PNP(Is=650.6E-18 Xti=3 Eg=1.11 Vaf=115.7 Bf=231.7 Ne=1.829 Ise=54.81f Ikf=1.079 Xtb=1.5 Br=3.563 Nc=2 Isc=0 Ikr=0 Rc=.715 Cjc=14.76p Mjc=.5383 Vjc=.75 Fc=.5 Cje=19.82p Mje=.3357 Vje=.75 Tr=111.3n Tf=603.7p Itf=.65 Vtf=5 Xtf=1.7 Rb=10 Vceo=60 Icrating=600m mfg=Philips)
.model 2N4401 NPN(Is=26.03f Xti=3 Eg=1.11 Vaf=90.7 Bf=4.292K Ne=1.244 Ise=26.03f Ikf=.2061 Xtb=1.5 Br=1.01 Nc=2 Isc=0 Ikr=0 Rc=.5 Cjc=11.01p Mjc=.3763 Vjc=.75 Fc=.5 Cje=24.07p Mje=.3641 Vje=.75 Tr=233.7n Tf=466.5p Itf=0 Vtf=0 Xtf=0 Rb=10 Vceo=40 Icrating=600m mfg=Fairchild)
.model 2N4403 PNP(Is=650.6E-18 Xti=3 Eg=1.11 Vaf=115.7 Bf=216.2 Ne=1.829 Ise=58.72f Ikf=1.079 Xtb=1.5 Br=3.578 Nc=2 Isc=0 Ikr=0 Rc=.715 Cjc=14.76p Mjc=.5383 Vjc=.75 Fc=.5 Cje=19.82p Mje=.3357 Vje=.75 Tr=111.6n Tf=603.7p Itf=.65 Vtf=5 Xtf=1.7 Rb=10 Vceo=40 Icrating=600m mfg=Fairchild)
.model 2N5550 NPN(Is=2.511f Xti=3 Eg=1.11 Vaf=100 Bf=213.4 Ne=1.241 Ise=2.511f Ikf=.3495 Xtb=1.5 Br=3.24 Nc=2 Isc=0 Ikr=0 Rc=1 Cjc=4.883p Mjc=.3047 Vjc=.75 Fc=.5 Cje=18.79p Mje=.3416 Vje=.75 Tr=1.212n Tf=560.1p Itf=50m Vtf=5 Xtf=8 Rb=10 Vceo=150 Icrating=600m mfg=Fairchild)
.model 2N5401 PNP(Is=21.48f Xti=3 Eg=1.11 Vaf=100 Bf=132.1 Ne=1.375 Ise=21.48f Ikf=.1848 Xtb=1.5 Br=3.661 Nc=2 Isc=0 Ikr=0 Rc=1.6 Cjc=17.63p Mjc=.5312 Vjc=.75 Fc=.5 Cje=73.39p Mje=.3777 Vje=.75 Tr=1.476n Tf=641.9p Itf=0 Vtf=0 Xtf=0 Rb=10 Vceo=150 Icrating=600m mfg=Fairchild)
.model 2N2369 NPN(Is=44.14f Xti=3 Eg=1.11 Vaf=100 Bf=78.32 Ne=1.389 Ise=91.95f Ikf=.3498 Xtb=1.5 Br=12.69m Nc=2 Isc=0 Ikr=0 Rc=.6 Cjc=2.83p Mjc=86.19m Vjc=.75 Fc=.5 Cje=4.5p Mje=.2418 Vje=.75 Tr=1.073u Tf=227.6p Itf=.3 Vtf=4 Xtf=4 Rb=10 Vceo=15 Icrating=200m mfg=Philips)
.model 2N5769 NPN(Is=44.14f Xti=3 Eg=1.11 Vaf=100 Bf=78.32 Ne=1.389 Ise=91.95f Ikf=.3498 Xtb=1.5 Br=12.69m Nc=2 Isc=0 Ikr=0 Rc=.6 Cjc=2.83p Mjc=86.19m Vjc=.75 Fc=.5 Cje=4.5p Mje=.2418 Vje=.75 Tr=1.073u Tf=227.6p Itf=.3 Vtf=4 Xtf=4 Rb=10 Vceo=15 Icrating=200m mfg=Fairchild)
.model 2N5771 PNP(Is=545.6E-18 Xti=3 Eg=1.11 Vaf=100 Bf=76.77 Ne=1.5 Ise=0 Ikf=50m Xtb=1.5 Br=1.365 Nc=2 Isc=0 Ikr=0 Rc=3.75 Cjc=2.77p Mjc=.1416 Vjc=.75 Fc=.5 Cje=2.65p Mje=.3083 Vje=.75 Tr=4.033n Tf=118.5p Itf=.5 Vtf=3 Xtf=6 Rb=10 Vceo=15 Icrating=200m mfg=Fairchild)
.model 2N3055 NPN(Bf=73 Br=2.66 Rb=.81 Rc=.0856 Re=.000856 CJC=1000P PC=.75 MC=.33 Tr=.5703U Is=2.37E-8 CJE=415P PE=.75 ME=.5 TF=99.52N NE=1.26 IK=1 Vceo=60 Icrating=10 mfg=STMicro)
.model BCW60A NPN(IS=20f VAF=100 BF=120 IKF=0.8 XTB=1.5 BR=5 CJC=20p CJE=8p TR=100n TF=600p RB=10 RC=3 RE=1 Vceo=32 Icrating=200m mfg=ROHM)
.model BCW60B NPN(IS=20f VAF=80 BF=240 IKF=1.0 XTB=1.5 BR=5 CJC=20p CJE=8p TR=100n TF=600p RB=10 RC=3 RE=1 Vceo=32 Icrating=200m mfg=ROHM)
.model BCW60C NPN(IS=20f VAF=65 BF=360 IKF=1.3 XTB=1.5 BR=5 CJC=20p CJE=8p TR=100n TF=600p RB=10 RC=3 RE=1 Vceo=32 Icrating=200m mfg=ROHM)
.model BCW60D NPN(IS=20f VAF=45 BF=500 IKF=1.5 XTB=1.5 BR=5 CJC=20p CJE=8p TR=100n TF=600p RB=10 RC=3 RE=1 Vceo=32 Icrating=200m mfg=ROHM)
.model BCW68F PNP(Is=40f VAF=100 Bf=175 IKF=2 Br=6 RC=.5 RE=0.1 RB=0.2 CJC=13p CJE=60p TR=12n TF=600p Vceo=45 Icrating=800m mfg=ROHM)
.model BCW68G PNP(Is=40f VAF=80 Bf=280 IKF=2.5 Br=6 RC=.5 RE=0.1 RB=0.2 CJC=13p CJE=60p TR=12n TF=600p Vceo=45 Icrating=800m mfg=ROHM)
.model BC547 NPN(Is=23.9f Xti=3 Eg=1.11 Vaf=63.2 Bf=294.3 Ne=1.541 Ise=3.545f Ikf=0.1357 Xtb=0 Br=7.946 Nc=1.243 Isc=62.72f Ikr=0.1144 Rc=0.85 Cjc=3.728p Mjc=.2955 Vjc=0.3997 Fc=.9579 Cje=13.58p Mje=0.3279 Vje=0.65 Tr=1E-32 Tf=0.4391n Itf=.7495 Vtf=2.643 Xtf=120 Rb=1 Nf=1.008 Nr=1.004 Var=25.9 Irb=1u Rbm=1 Re=0.4683 Cjs=0 Vjs=0.75 Mjs=0.333 Vceo=45 Icrating=100m mfg=Philips)
.model BC557 PNP(Is=38.34f Xti=3 Eg=1.11 Vaf=21.11 Bf=344.4 Ne=1.528 Ise=12.19f Ikf=0.08039 Xtb=0 Br=14.84 Nc=1.28 Isc=285.2f Ikr=0.047 Rc=0.5713 Cjc=10.84p Mjc=.3563 Vjc=0.1022 Fc=.8027 Cje=12.3p Mje=0.378 Vje=0.6016 Tr=1E-32 Tf=0.5595n Itf=0.1483 Vtf=5.23 Xtf=3.414 Rb=1 Nf=1.008 Nr=1.005 Var=32.02 Irb=1u Rbm=1 Re=0.6202 Cjs=0 Vjs=0.75 Mjs=0.333 Vceo=45 Icrating=100m mfg=Philips)
.model MJF15030 NPN(Is=8.52586e-11 Bf=111.756 Nf=1.12559 Vaf=24.6951 Ikf=9.20535 Ise=5.49997e-12 Ne=3.4375 Br=3.01415 Nr=1.24186 Var=3.47825 Ikr=6.10635 Isc=6.25e-13 Nc=3.90625 Rb=8.46485 Irb=0.1 Rbm=0.1 Re=0.00048424 Rc=0.142581 Xtb=0.120563 Xti=1 Eg=1.10791 Cje=3.00414e-09 Vje=0.411662 Mje=0.51835 Tf=1.87342e-09 Xtf=1000 Vtf=2395.66 Itf=178.85 Cjc=2.59252e-10 Vjc=0.4 Mjc=0.383014 Xcjc=0.785372 Fc=0.1 Cjs=0 Vjs=0.75 Mjs=0.5 Tr=8.8568e-07 Ptf=0 Kf=0 Af=1 Vceo=150 Icrating=8)
.model MJF15031 PNP(Is=8.44385e-11,bf=118.835,nf=1.22766,vaf=24.5822,ikf=9.15247,ise=5.49989e-12,ne=3.43751,br=2.98261,nr=1.41393,var=3.42026,ikr=6.68823,isc=6.25e-13,nc=3.90625,rb=8.19612,irb=0.1,rbm=0.1,re=0.000474198,rc=0.125756,xtb=0.120732,xti=1,eg=1.10974,cje=1.55377e-09,vje=0.99,mje=0.547635,tf=6.50306e-10,xtf=30.1354,vtf=2.33133,itf=0.0183389,cjc=5e-10,vjc=0.4,mjc=0.411581,xcjc=0.793472,fc=0.1,cjs=0,vjs=0.75,mjs=0.5,tr=7.75795e-07,ptf=0,kf=0,af=1 Vceo=150 Icrating=8)
.model CA3086 NPN(Is=10f Xti=3 Eg=1.11 Vaf=100 VAR=1.000E + 02 Bf=156.6 Ise=114.886f Ne=1.47 Ikf=36.7M Xtb=0.0 Br=.1 Isc=10f Nc=2 Ikr=10M Rc=10 Cjc=991.79f Mjc=0.333 Vjc=0.75 Fc=0.5 Cje=1.02p Mje=.336 Vje=0.75 Tr=10n Tf=278.55n Itf=.77 Xtf=91.38 Vtf=18.37 Ptf=0 Re=0 Rb=0)
.MODEL QBC558A/PLP PNP(IS=20.59f NF=1.003 ISE=2.971E-15 NE=1.316 BF=227.3 IKF=0.08719 VAF=37.2 NR=1.007 ISC=1.339E-14 NC=1.15 BR=7.69 IKR=0.07646 VAR=11.42 RB=1 IRB=1E-06 RBM=1 RE=0.688 RC=0.6437 XTB=0 EG=1.11 XTI=3 CJE=1.4E-11 VJE=0.5912 MJE=0.3572 TF=7.046E-10 XTF=4.217 VTF=5.367 ITF=0.1947 PTF=0 CJC=1.113E-11 VJC=0.1 MJC=0.3414 XCJC=0.6288 TR=1E-32 CJS=0 VJS=0.75 MJS=0.333 FC=0.7947 Vceo=30 Icrating=100m)
.MODEL QBC548B/PLP NPN(IS=23.9f NF=1.008 ISE=3.545E-15 NE=1.541 BF=294.3 IKF=0.1357 VAF=63.2 NR=1.004 ISC=6.272E-14 NC=1.243 BR=7.946 IKR=0.1144 VAR=25.9 RB=1 IRB=1E-06 RBM=1 RE=0.4683 RC=0.85 XTB=0 EG=1.11 XTI=3 CJE=1.358E-11 VJE=0.65 MJE=0.3279 TF=4.391E-10 XTF=120 VTF=2.643 ITF=0.7495 PTF=0 CJC=3.728E-12 VJC=0.3997 MJC=0.2955 XCJC=0.6193 TR=1E-32 CJS=0 VJS=0.75 MJS=0.333 FC=0.9579 Vceo=30 Icrating=100m)
.MODEL QBD139 npn(IS=1e-09 BF=222.664 NF=0.85 VAF=36.4079 IKF=0.166126 ISE=5.03418e-09 NE=1.45313 BR=1.35467 NR=1.33751 VAR=142.931 IKR=1.66126 ISC=5.02557e-09 NC=3.10227 RB=26.9143 IRB=0.1 RBM=0.1 RE=0.000472454 RC=1.04109 XTB=0.727762 XTI=1.04311 EG=1.05 CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09 XTF=1 VTF=10 ITF=0.01 CJC=1e-11 VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1 Vceo=80 Icrating=1000m)
.model 2N3019 NPN(Is=14f Vaf=100 Bf=200 Ikf=.75 Xtb=1.5 Br=5 Rc=.7 Cjc=16p Mjc=.36 Cje=55p Mje=.1553 Tr=800p Tf=800p Itf=1.2 Vtf=5 Xtf=55 Rb=10 Vceo=80 Icrating=1 mfg=Semicoa)
.MODEL QBD140 pnp(IS=1e-09 BF=650.842 NF=0.85 VAF=10 IKF=0.0950125 ISE=1e-08 NE=1.54571 BR=56.177 NR=1.5 VAR=2.11267 IKR=0.950125 ISC=1e-08 NC=3.58527 RB=41.7566 IRB=0.1 RBM=0.108893 RE=0.000347052 RC=1.32566 XTB=19.5239 XTI=1 EG=1.05 CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09 XTF=1 VTF=10 ITF=0.01CJC=1e-11 VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1 Vceo=80 Icrating=1000m)
.MODEL QMJE3055t npn(IS=1.92238e-13 BF=327.43 NF=0.85 VAF=36.105 IKF=0.620037 ISE=1.4602e-10 NE=1.50926 BR=0.654697 NR=0.935367 VAR=361.05 IKR=6.20037 ISC=6.85154e-12 NC=2.96871 RB=16.05 IRB=0.1 RBM=0.161446 RE=0.000602331 RC=0.0632768 XTB=0.943656 XTI=1.12302 EG=1.05 CJE=9.23675e-08 VJE=0.506151 MJE=0.607139 TF=1e-08 XTF=1.35736 VTF=0.997047 ITF=0.999796 CJC=5e-10 VJC=0.400198 MJC=0.410184 XCJC=0.803125 FC=0.658133 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1)
.MODEL QMJE2955t pnp(IS=4.14254e-10 BF=449.16 NF=0.85 VAF=17.4911 IKF=0.414206 ISE=1e-08 NE=1.47014 BR=0.1 NR=1.09325 VAR=174.911 IKR=4.14206 ISC=7.59792e-09 NC=3.02799 RB=20.1795 IRB=0.1 RBM=0.1 RE=0.000499379 RC=0.0813684 XTB=0.1 XTI=1.16399 EG=1.05 CJE=9.97416e-08 VJE=0.416937 MJE=0.61618 TF=9.98874e-09 XTF=1.35736 VTF=0.997021 ITF=0.999788 CJC=4.99998e-10 VJC=0.40025 MJC=0.410011 XCJC=0.803124 FC=0.661649 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1)
.MODEL Qtip31 npn (IS=1e-09 BF=3656.16 NF=1.23899 VAF=10 IKF=0.0333653 ISE=1e-08 NE=2.29374 BR=0.1 NR=1.5 VAR=100 IKR=0.333653 ISC=1e-08 NC=1.75728 RB=6.15083 IRB=100 RBM=0.00113049 RE=0.0001 RC=0.0491489 XTB=50 XTI=1 EG=1.05 CJE=3.26475e-10 VJE=0.446174 MJE=0.464221 TF=2.06218e-09 XTF=15.0842 VTF=25.7317 ITF=0.001 CJC=3.07593e-10 VJC=0.775484 MJC=0.476498 XCJC=0.750493 FC=0.796407 CJS=0 VJS=0.75 MJS=0.5 TR=9.57121e-06 PTF=0 KF=0 AF=1)
.MODEL Qtip32c pnp (IS=1e-09 BF=134.366 NF=1.29961 VAF=10 IKF=0.742988 ISE=1e-16 NE=1.40014 BR=0.1 NR=1.46599 VAR=100 IKR=3.21978 ISC=1e-16 NC=2.71657 RB=7.44433 IRB=2.41268 RBM=0.218936 RE=0.0152284 RC=0.0761421 XTB=0.1 XTI=1 EG=1.05 CJE=3.26474e-10 VJE=0.446178 MJE=0.464223 TF=1e-08 XTF=3.50642 VTF=8.2848 ITF=0.0305862 CJC=3.07595e-10 VJC=0.77548 MJC=0.476497 XCJC=0.799334 FC=0.8 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1)
.MODEL q2n3906 pnp (IS=7.75521e-12 BF=194.093 NF=1.35509 VAF=156.436 IKF=0.0660057 ISE=1.88546e-12 NE=1.81673 BR=3.41317 NR=1.5 VAR=5.86061 IKR=1.70599 ISC=7.64281e-10 NC=1.92376 RB=6.48961 IRB=0.1 RBM=0.1 RE=0.0001 RC=2.45044 XTB=0.1 XTI=1 EG=1.05 CJE=6.11928e-12 VJE=0.4 MJE=0.248812 TF=5.21843e-10 XTF=0.932702 VTF=9.1046 ITF=0.0106472 CJC=6.85007e-12 VJC=0.4 MJC=0.279018 XCJC=0.9 FC=0.478887 CJS=0 VJS=0.75 MJS=0.5 TR=4.30605e-07 PTF=0 KF=0 AF=1)

* hello
